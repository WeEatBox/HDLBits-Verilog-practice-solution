module top_module( input in, output out );
    not n1(out,in); // build-in not gate module
endmodule