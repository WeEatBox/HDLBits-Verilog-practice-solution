module top_module (
    input [3:0] SW,
    input [3:0] KEY,
    output [3:0] LEDR
); //

    MUXDFF m_0(KEY[0],LEDR[1],SW[0],KEY[1],KEY[2],LEDR[0]);
    MUXDFF m_1(KEY[0],LEDR[2],SW[1],KEY[1],KEY[2],LEDR[1]);
    MUXDFF m_2(KEY[0],LEDR[3],SW[2],KEY[1],KEY[2],LEDR[2]);
    MUXDFF m_3(KEY[0],KEY[3],SW[3],KEY[1],KEY[2],LEDR[3]);
  
endmodule

module MUXDFF (
    input clk,
    input w, R, E, L,
    output Q
);
    wire tmp0,tmp1;
    assign tmp0 = E? w: Q;
    assign tmp1 = L? R: tmp0;
    
    always@(posedge clk) Q <= tmp1;
endmodule
